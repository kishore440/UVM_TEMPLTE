module tb;
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "uvm_pkg.sv"
initial
begin
        run_test("my_test");
end
endmodule
